`ifndef SPI_DEFINE
`define SPI_DEFINE

`define BIT_ADDR_NUM 4
`define BIT_DATA_NUM 8
`define BIT_FULL_SIZE 16

`endif